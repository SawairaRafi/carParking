library verilog;
use verilog.vl_types.all;
entity car_parking_system_vlg_vec_tst is
end car_parking_system_vlg_vec_tst;
